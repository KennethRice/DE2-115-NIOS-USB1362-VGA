// DE2_115_SOPC.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module DE2_115_SOPC (
		output wire        altpll_sys,                   //               c0_out_clk.clk
		output wire        altpll_io,                    //               c2_out_clk.clk
		output wire        c3_out_clk_clk,               //               c3_out_clk.clk
		input  wire        clk_50,                       //            clk_50_clk_in.clk
		input  wire        reset_n,                      //      clk_50_clk_in_reset.reset_n
		input  wire [3:0]  in_port_to_the_key,           //  key_external_connection.export
		output wire        LCD_RS_from_the_lcd,          //             lcd_external.RS
		output wire        LCD_RW_from_the_lcd,          //                         .RW
		inout  wire [7:0]  LCD_data_to_and_from_the_lcd, //                         .data
		output wire        LCD_E_from_the_lcd,           //                         .E
		output wire [8:0]  out_port_from_the_ledg,       // ledg_external_connection.export
		output wire [17:0] out_port_from_the_ledr,       // ledr_external_connection.export
		input  wire        pll_areset_conduit_export,    //       pll_areset_conduit.export
		output wire        altpll_sdram,                 //                   pll_c1.clk
		output wire        locked_from_the_pll,          //       pll_locked_conduit.export
		output wire [12:0] zs_addr_from_the_sdram,       //               sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,         //                         .ba
		output wire        zs_cas_n_from_the_sdram,      //                         .cas_n
		output wire        zs_cke_from_the_sdram,        //                         .cke
		output wire        zs_cs_n_from_the_sdram,       //                         .cs_n
		inout  wire [31:0] zs_dq_to_and_from_the_sdram,  //                         .dq
		output wire [3:0]  zs_dqm_from_the_sdram,        //                         .dqm
		output wire        zs_ras_n_from_the_sdram,      //                         .ras_n
		output wire        zs_we_n_from_the_sdram,       //                         .we_n
		output wire [63:0] SEG7_from_the_seg7,           //         seg7_conduit_end.export
		input  wire [17:0] in_port_to_the_sw,            //   sw_external_connection.export
		inout  wire [15:0] usb_conduit_end_DATA,         //          usb_conduit_end.DATA
		output wire [1:0]  usb_conduit_end_ADDR,         //                         .ADDR
		output wire        usb_conduit_end_RD_N,         //                         .RD_N
		output wire        usb_conduit_end_WR_N,         //                         .WR_N
		output wire        usb_conduit_end_CS_N,         //                         .CS_N
		output wire        usb_conduit_end_RST_N,        //                         .RST_N
		input  wire        usb_conduit_end_INT0,         //                         .INT0
		input  wire        usb_conduit_end_INT1,         //                         .INT1
		output wire        vga_data_CLK,                 //                 vga_data.CLK
		output wire        vga_data_HS,                  //                         .HS
		output wire        vga_data_VS,                  //                         .VS
		output wire        vga_data_BLANK,               //                         .BLANK
		output wire        vga_data_SYNC,                //                         .SYNC
		output wire [7:0]  vga_data_R,                   //                         .R
		output wire [7:0]  vga_data_G,                   //                         .G
		output wire [7:0]  vga_data_B                    //                         .B
	);

	wire         video_rgb_resampler_0_avalon_rgb_source_valid;             // video_rgb_resampler_0:stream_out_valid -> vga:valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;              // video_rgb_resampler_0:stream_out_data -> vga:data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;             // vga:ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;     // video_rgb_resampler_0:stream_out_startofpacket -> vga:startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;       // video_rgb_resampler_0:stream_out_endofpacket -> vga:endofpacket
	wire         lcd_ta_sgdma_to_fifo_out_valid;                            // lcd_ta_sgdma_to_fifo:out_valid -> lcd_pixel_fifo:avalonst_sink_valid
	wire  [63:0] lcd_ta_sgdma_to_fifo_out_data;                             // lcd_ta_sgdma_to_fifo:out_data -> lcd_pixel_fifo:avalonst_sink_data
	wire         lcd_ta_sgdma_to_fifo_out_ready;                            // lcd_pixel_fifo:avalonst_sink_ready -> lcd_ta_sgdma_to_fifo:out_ready
	wire         lcd_ta_sgdma_to_fifo_out_startofpacket;                    // lcd_ta_sgdma_to_fifo:out_startofpacket -> lcd_pixel_fifo:avalonst_sink_startofpacket
	wire         lcd_ta_sgdma_to_fifo_out_endofpacket;                      // lcd_ta_sgdma_to_fifo:out_endofpacket -> lcd_pixel_fifo:avalonst_sink_endofpacket
	wire   [2:0] lcd_ta_sgdma_to_fifo_out_empty;                            // lcd_ta_sgdma_to_fifo:out_empty -> lcd_pixel_fifo:avalonst_sink_empty
	wire         lcd_pixel_fifo_out_valid;                                  // lcd_pixel_fifo:avalonst_source_valid -> lcd_ta_fifo_to_dfa:in_valid
	wire  [63:0] lcd_pixel_fifo_out_data;                                   // lcd_pixel_fifo:avalonst_source_data -> lcd_ta_fifo_to_dfa:in_data
	wire         lcd_pixel_fifo_out_ready;                                  // lcd_ta_fifo_to_dfa:in_ready -> lcd_pixel_fifo:avalonst_source_ready
	wire         lcd_pixel_fifo_out_startofpacket;                          // lcd_pixel_fifo:avalonst_source_startofpacket -> lcd_ta_fifo_to_dfa:in_startofpacket
	wire         lcd_pixel_fifo_out_endofpacket;                            // lcd_pixel_fifo:avalonst_source_endofpacket -> lcd_ta_fifo_to_dfa:in_endofpacket
	wire   [2:0] lcd_pixel_fifo_out_empty;                                  // lcd_pixel_fifo:avalonst_source_empty -> lcd_ta_fifo_to_dfa:in_empty
	wire         lcd_ta_fifo_to_dfa_out_valid;                              // lcd_ta_fifo_to_dfa:out_valid -> lcd_64_to_8_bits_dfa:in_valid
	wire  [63:0] lcd_ta_fifo_to_dfa_out_data;                               // lcd_ta_fifo_to_dfa:out_data -> lcd_64_to_8_bits_dfa:in_data
	wire         lcd_ta_fifo_to_dfa_out_ready;                              // lcd_64_to_8_bits_dfa:in_ready -> lcd_ta_fifo_to_dfa:out_ready
	wire         lcd_ta_fifo_to_dfa_out_startofpacket;                      // lcd_ta_fifo_to_dfa:out_startofpacket -> lcd_64_to_8_bits_dfa:in_startofpacket
	wire         lcd_ta_fifo_to_dfa_out_endofpacket;                        // lcd_ta_fifo_to_dfa:out_endofpacket -> lcd_64_to_8_bits_dfa:in_endofpacket
	wire   [2:0] lcd_ta_fifo_to_dfa_out_empty;                              // lcd_ta_fifo_to_dfa:out_empty -> lcd_64_to_8_bits_dfa:in_empty
	wire         lcd_64_to_8_bits_dfa_out_valid;                            // lcd_64_to_8_bits_dfa:out_valid -> lcd_pixel_converter:valid_in
	wire  [31:0] lcd_64_to_8_bits_dfa_out_data;                             // lcd_64_to_8_bits_dfa:out_data -> lcd_pixel_converter:data_in
	wire         lcd_64_to_8_bits_dfa_out_ready;                            // lcd_pixel_converter:ready_out -> lcd_64_to_8_bits_dfa:out_ready
	wire         lcd_64_to_8_bits_dfa_out_startofpacket;                    // lcd_64_to_8_bits_dfa:out_startofpacket -> lcd_pixel_converter:sop_in
	wire         lcd_64_to_8_bits_dfa_out_endofpacket;                      // lcd_64_to_8_bits_dfa:out_endofpacket -> lcd_pixel_converter:eop_in
	wire   [1:0] lcd_64_to_8_bits_dfa_out_empty;                            // lcd_64_to_8_bits_dfa:out_empty -> lcd_pixel_converter:empty_in
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] lcd_sgdma_descriptor_read_readdata;                        // mm_interconnect_0:lcd_sgdma_descriptor_read_readdata -> lcd_sgdma:descriptor_read_readdata
	wire         lcd_sgdma_descriptor_read_waitrequest;                     // mm_interconnect_0:lcd_sgdma_descriptor_read_waitrequest -> lcd_sgdma:descriptor_read_waitrequest
	wire  [31:0] lcd_sgdma_descriptor_read_address;                         // lcd_sgdma:descriptor_read_address -> mm_interconnect_0:lcd_sgdma_descriptor_read_address
	wire         lcd_sgdma_descriptor_read_read;                            // lcd_sgdma:descriptor_read_read -> mm_interconnect_0:lcd_sgdma_descriptor_read_read
	wire         lcd_sgdma_descriptor_read_readdatavalid;                   // mm_interconnect_0:lcd_sgdma_descriptor_read_readdatavalid -> lcd_sgdma:descriptor_read_readdatavalid
	wire         lcd_sgdma_descriptor_write_waitrequest;                    // mm_interconnect_0:lcd_sgdma_descriptor_write_waitrequest -> lcd_sgdma:descriptor_write_waitrequest
	wire  [31:0] lcd_sgdma_descriptor_write_address;                        // lcd_sgdma:descriptor_write_address -> mm_interconnect_0:lcd_sgdma_descriptor_write_address
	wire         lcd_sgdma_descriptor_write_write;                          // lcd_sgdma:descriptor_write_write -> mm_interconnect_0:lcd_sgdma_descriptor_write_write
	wire  [31:0] lcd_sgdma_descriptor_write_writedata;                      // lcd_sgdma:descriptor_write_writedata -> mm_interconnect_0:lcd_sgdma_descriptor_write_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] lcd_sgdma_m_read_readdata;                                 // mm_interconnect_0:lcd_sgdma_m_read_readdata -> lcd_sgdma:m_read_readdata
	wire         lcd_sgdma_m_read_waitrequest;                              // mm_interconnect_0:lcd_sgdma_m_read_waitrequest -> lcd_sgdma:m_read_waitrequest
	wire  [31:0] lcd_sgdma_m_read_address;                                  // lcd_sgdma:m_read_address -> mm_interconnect_0:lcd_sgdma_m_read_address
	wire         lcd_sgdma_m_read_read;                                     // lcd_sgdma:m_read_read -> mm_interconnect_0:lcd_sgdma_m_read_read
	wire         lcd_sgdma_m_read_readdatavalid;                            // mm_interconnect_0:lcd_sgdma_m_read_readdatavalid -> lcd_sgdma:m_read_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_lcd_sgdma_csr_chipselect;                // mm_interconnect_0:lcd_sgdma_csr_chipselect -> lcd_sgdma:csr_chipselect
	wire  [31:0] mm_interconnect_0_lcd_sgdma_csr_readdata;                  // lcd_sgdma:csr_readdata -> mm_interconnect_0:lcd_sgdma_csr_readdata
	wire   [3:0] mm_interconnect_0_lcd_sgdma_csr_address;                   // mm_interconnect_0:lcd_sgdma_csr_address -> lcd_sgdma:csr_address
	wire         mm_interconnect_0_lcd_sgdma_csr_read;                      // mm_interconnect_0:lcd_sgdma_csr_read -> lcd_sgdma:csr_read
	wire         mm_interconnect_0_lcd_sgdma_csr_write;                     // mm_interconnect_0:lcd_sgdma_csr_write -> lcd_sgdma:csr_write
	wire  [31:0] mm_interconnect_0_lcd_sgdma_csr_writedata;                 // mm_interconnect_0:lcd_sgdma_csr_writedata -> lcd_sgdma:csr_writedata
	wire         mm_interconnect_0_isp1362_if_0_dc_chipselect;              // mm_interconnect_0:ISP1362_IF_0_dc_chipselect -> ISP1362_IF_0:avs_dc_chipselect_n_iCS_N
	wire  [15:0] mm_interconnect_0_isp1362_if_0_dc_readdata;                // ISP1362_IF_0:avs_dc_readdata_oDATA -> mm_interconnect_0:ISP1362_IF_0_dc_readdata
	wire   [0:0] mm_interconnect_0_isp1362_if_0_dc_address;                 // mm_interconnect_0:ISP1362_IF_0_dc_address -> ISP1362_IF_0:avs_dc_address_iADDR
	wire         mm_interconnect_0_isp1362_if_0_dc_read;                    // mm_interconnect_0:ISP1362_IF_0_dc_read -> ISP1362_IF_0:avs_dc_read_n_iRD_N
	wire         mm_interconnect_0_isp1362_if_0_dc_write;                   // mm_interconnect_0:ISP1362_IF_0_dc_write -> ISP1362_IF_0:avs_dc_write_n_iWR_N
	wire  [15:0] mm_interconnect_0_isp1362_if_0_dc_writedata;               // mm_interconnect_0:ISP1362_IF_0_dc_writedata -> ISP1362_IF_0:avs_dc_writedata_iDATA
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_isp1362_if_0_hc_chipselect;              // mm_interconnect_0:ISP1362_IF_0_hc_chipselect -> ISP1362_IF_0:avs_hc_chipselect_n_iCS_N
	wire  [15:0] mm_interconnect_0_isp1362_if_0_hc_readdata;                // ISP1362_IF_0:avs_hc_readdata_oDATA -> mm_interconnect_0:ISP1362_IF_0_hc_readdata
	wire   [0:0] mm_interconnect_0_isp1362_if_0_hc_address;                 // mm_interconnect_0:ISP1362_IF_0_hc_address -> ISP1362_IF_0:avs_hc_address_iADDR
	wire         mm_interconnect_0_isp1362_if_0_hc_read;                    // mm_interconnect_0:ISP1362_IF_0_hc_read -> ISP1362_IF_0:avs_hc_read_n_iRD_N
	wire         mm_interconnect_0_isp1362_if_0_hc_write;                   // mm_interconnect_0:ISP1362_IF_0_hc_write -> ISP1362_IF_0:avs_hc_write_n_iWR_N
	wire  [15:0] mm_interconnect_0_isp1362_if_0_hc_writedata;               // mm_interconnect_0:ISP1362_IF_0_hc_writedata -> ISP1362_IF_0:avs_hc_writedata_iDATA
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                  // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                   // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                      // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                     // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                 // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_readdata;           // clock_crossing_io:s0_readdata -> mm_interconnect_0:clock_crossing_io_s0_readdata
	wire         mm_interconnect_0_clock_crossing_io_s0_waitrequest;        // clock_crossing_io:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_s0_waitrequest
	wire         mm_interconnect_0_clock_crossing_io_s0_debugaccess;        // mm_interconnect_0:clock_crossing_io_s0_debugaccess -> clock_crossing_io:s0_debugaccess
	wire  [21:0] mm_interconnect_0_clock_crossing_io_s0_address;            // mm_interconnect_0:clock_crossing_io_s0_address -> clock_crossing_io:s0_address
	wire         mm_interconnect_0_clock_crossing_io_s0_read;               // mm_interconnect_0:clock_crossing_io_s0_read -> clock_crossing_io:s0_read
	wire   [3:0] mm_interconnect_0_clock_crossing_io_s0_byteenable;         // mm_interconnect_0:clock_crossing_io_s0_byteenable -> clock_crossing_io:s0_byteenable
	wire         mm_interconnect_0_clock_crossing_io_s0_readdatavalid;      // clock_crossing_io:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_s0_readdatavalid
	wire         mm_interconnect_0_clock_crossing_io_s0_write;              // mm_interconnect_0:clock_crossing_io_s0_write -> clock_crossing_io:s0_write
	wire  [31:0] mm_interconnect_0_clock_crossing_io_s0_writedata;          // mm_interconnect_0:clock_crossing_io_s0_writedata -> clock_crossing_io:s0_writedata
	wire   [0:0] mm_interconnect_0_clock_crossing_io_s0_burstcount;         // mm_interconnect_0:clock_crossing_io_s0_burstcount -> clock_crossing_io:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_stamp_s1_chipselect;               // mm_interconnect_0:timer_stamp_s1_chipselect -> timer_stamp:chipselect
	wire  [15:0] mm_interconnect_0_timer_stamp_s1_readdata;                 // timer_stamp:readdata -> mm_interconnect_0:timer_stamp_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_stamp_s1_address;                  // mm_interconnect_0:timer_stamp_s1_address -> timer_stamp:address
	wire         mm_interconnect_0_timer_stamp_s1_write;                    // mm_interconnect_0:timer_stamp_s1_write -> timer_stamp:write_n
	wire  [15:0] mm_interconnect_0_timer_stamp_s1_writedata;                // mm_interconnect_0:timer_stamp_s1_writedata -> timer_stamp:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         clock_crossing_io_m0_waitrequest;                          // mm_interconnect_1:clock_crossing_io_m0_waitrequest -> clock_crossing_io:m0_waitrequest
	wire  [31:0] clock_crossing_io_m0_readdata;                             // mm_interconnect_1:clock_crossing_io_m0_readdata -> clock_crossing_io:m0_readdata
	wire         clock_crossing_io_m0_debugaccess;                          // clock_crossing_io:m0_debugaccess -> mm_interconnect_1:clock_crossing_io_m0_debugaccess
	wire  [21:0] clock_crossing_io_m0_address;                              // clock_crossing_io:m0_address -> mm_interconnect_1:clock_crossing_io_m0_address
	wire         clock_crossing_io_m0_read;                                 // clock_crossing_io:m0_read -> mm_interconnect_1:clock_crossing_io_m0_read
	wire   [3:0] clock_crossing_io_m0_byteenable;                           // clock_crossing_io:m0_byteenable -> mm_interconnect_1:clock_crossing_io_m0_byteenable
	wire         clock_crossing_io_m0_readdatavalid;                        // mm_interconnect_1:clock_crossing_io_m0_readdatavalid -> clock_crossing_io:m0_readdatavalid
	wire  [31:0] clock_crossing_io_m0_writedata;                            // clock_crossing_io:m0_writedata -> mm_interconnect_1:clock_crossing_io_m0_writedata
	wire         clock_crossing_io_m0_write;                                // clock_crossing_io:m0_write -> mm_interconnect_1:clock_crossing_io_m0_write
	wire   [0:0] clock_crossing_io_m0_burstcount;                           // clock_crossing_io:m0_burstcount -> mm_interconnect_1:clock_crossing_io_m0_burstcount
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_readdata;              // seg7:s_readdata -> mm_interconnect_1:seg7_avalon_slave_readdata
	wire   [2:0] mm_interconnect_1_seg7_avalon_slave_address;               // mm_interconnect_1:seg7_avalon_slave_address -> seg7:s_address
	wire         mm_interconnect_1_seg7_avalon_slave_read;                  // mm_interconnect_1:seg7_avalon_slave_read -> seg7:s_read
	wire         mm_interconnect_1_seg7_avalon_slave_write;                 // mm_interconnect_1:seg7_avalon_slave_write -> seg7:s_write
	wire   [7:0] mm_interconnect_1_seg7_avalon_slave_writedata;             // mm_interconnect_1:seg7_avalon_slave_writedata -> seg7:s_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;             // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire   [7:0] mm_interconnect_1_lcd_control_slave_readdata;              // lcd:readdata -> mm_interconnect_1:lcd_control_slave_readdata
	wire   [1:0] mm_interconnect_1_lcd_control_slave_address;               // mm_interconnect_1:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_1_lcd_control_slave_read;                  // mm_interconnect_1:lcd_control_slave_read -> lcd:read
	wire         mm_interconnect_1_lcd_control_slave_begintransfer;         // mm_interconnect_1:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         mm_interconnect_1_lcd_control_slave_write;                 // mm_interconnect_1:lcd_control_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_1_lcd_control_slave_writedata;             // mm_interconnect_1:lcd_control_slave_writedata -> lcd:writedata
	wire         mm_interconnect_1_key_s1_chipselect;                       // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                         // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                          // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_write;                            // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                        // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire         mm_interconnect_1_sw_s1_chipselect;                        // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                          // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                           // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_write;                             // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                         // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_1_ledg_s1_chipselect;                      // mm_interconnect_1:ledg_s1_chipselect -> ledg:chipselect
	wire  [31:0] mm_interconnect_1_ledg_s1_readdata;                        // ledg:readdata -> mm_interconnect_1:ledg_s1_readdata
	wire   [1:0] mm_interconnect_1_ledg_s1_address;                         // mm_interconnect_1:ledg_s1_address -> ledg:address
	wire         mm_interconnect_1_ledg_s1_write;                           // mm_interconnect_1:ledg_s1_write -> ledg:write_n
	wire  [31:0] mm_interconnect_1_ledg_s1_writedata;                       // mm_interconnect_1:ledg_s1_writedata -> ledg:writedata
	wire         mm_interconnect_1_ledr_s1_chipselect;                      // mm_interconnect_1:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_1_ledr_s1_readdata;                        // ledr:readdata -> mm_interconnect_1:ledr_s1_readdata
	wire   [1:0] mm_interconnect_1_ledr_s1_address;                         // mm_interconnect_1:ledr_s1_address -> ledr:address
	wire         mm_interconnect_1_ledr_s1_write;                           // mm_interconnect_1:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_1_ledr_s1_writedata;                       // mm_interconnect_1:ledr_s1_writedata -> ledr:writedata
	wire         irq_mapper_receiver0_irq;                                  // lcd_sgdma:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // ISP1362_IF_0:avs_dc_irq_n_oINT0_N -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // ISP1362_IF_0:avs_hc_irq_n_oINT0_N -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver6_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                  // timer_stamp:irq -> irq_mapper:receiver7_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         irq_mapper_receiver3_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // timer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver4_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                         // key:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver5_irq;                                  // irq_synchronizer_002:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                         // sw:irq -> irq_synchronizer_002:receiver_irq
	wire         lcd_pixel_converter_out_valid;                             // lcd_pixel_converter:valid_out -> avalon_st_adapter:in_0_valid
	wire  [23:0] lcd_pixel_converter_out_data;                              // lcd_pixel_converter:data_out -> avalon_st_adapter:in_0_data
	wire         lcd_pixel_converter_out_ready;                             // avalon_st_adapter:in_0_ready -> lcd_pixel_converter:ready_in
	wire         lcd_pixel_converter_out_startofpacket;                     // lcd_pixel_converter:sop_out -> avalon_st_adapter:in_0_startofpacket
	wire         lcd_pixel_converter_out_endofpacket;                       // lcd_pixel_converter:eop_out -> avalon_st_adapter:in_0_endofpacket
	wire   [1:0] lcd_pixel_converter_out_empty;                             // lcd_pixel_converter:empty_out -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                             // avalon_st_adapter:out_0_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [23:0] avalon_st_adapter_out_0_data;                              // avalon_st_adapter:out_0_data -> video_rgb_resampler_0:stream_in_data
	wire         avalon_st_adapter_out_0_ready;                             // video_rgb_resampler_0:stream_in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                     // avalon_st_adapter:out_0_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                       // avalon_st_adapter:out_0_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         lcd_sgdma_out_valid;                                       // lcd_sgdma:out_valid -> avalon_st_adapter_001:in_0_valid
	wire  [31:0] lcd_sgdma_out_data;                                        // lcd_sgdma:out_data -> avalon_st_adapter_001:in_0_data
	wire         lcd_sgdma_out_ready;                                       // avalon_st_adapter_001:in_0_ready -> lcd_sgdma:out_ready
	wire         lcd_sgdma_out_startofpacket;                               // lcd_sgdma:out_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire         lcd_sgdma_out_endofpacket;                                 // lcd_sgdma:out_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire   [1:0] lcd_sgdma_out_empty;                                       // lcd_sgdma:out_empty -> avalon_st_adapter_001:in_0_empty
	wire         avalon_st_adapter_001_out_0_valid;                         // avalon_st_adapter_001:out_0_valid -> lcd_ta_sgdma_to_fifo:in_valid
	wire  [63:0] avalon_st_adapter_001_out_0_data;                          // avalon_st_adapter_001:out_0_data -> lcd_ta_sgdma_to_fifo:in_data
	wire         avalon_st_adapter_001_out_0_ready;                         // lcd_ta_sgdma_to_fifo:in_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;                 // avalon_st_adapter_001:out_0_startofpacket -> lcd_ta_sgdma_to_fifo:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;                   // avalon_st_adapter_001:out_0_endofpacket -> lcd_ta_sgdma_to_fifo:in_endofpacket
	wire   [2:0] avalon_st_adapter_001_out_0_empty;                         // avalon_st_adapter_001:out_0_empty -> lcd_ta_sgdma_to_fifo:in_empty
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [ISP1362_IF_0:avs_dc_reset_n_iRST_N, ISP1362_IF_0:avs_hc_reset_n_iRST_N, avalon_st_adapter_001:in_rst_0_reset, clock_crossing_io:s0_reset, cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, jtag_uart:rst_n, lcd_pixel_fifo:wrreset_n, lcd_sgdma:system_reset_n, lcd_ta_sgdma_to_fifo:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, timer_stamp:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [clock_crossing_io:m0_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, key:reset_n, lcd:reset_n, ledg:reset_n, ledr:reset_n, mm_interconnect_0:timer_reset_reset_bridge_in_reset_reset, mm_interconnect_1:clock_crossing_io_m0_reset_reset_bridge_in_reset_reset, seg7:s_reset, sw:reset_n, sysid:reset_n, timer:reset_n]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [avalon_st_adapter:in_rst_0_reset, lcd_64_to_8_bits_dfa:reset_n, lcd_pixel_converter:reset_n, lcd_pixel_fifo:rdreset_n, lcd_ta_fifo_to_dfa:reset_n, vga:reset, video_rgb_resampler_0:reset]
	wire         rst_controller_003_reset_out_reset;                        // rst_controller_003:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	ISP1362_IF isp1362_if_0 (
		.avs_hc_clk_iCLK           (altpll_sys),                                    //       hc_clock.clk
		.avs_hc_reset_n_iRST_N     (~rst_controller_reset_out_reset),               // hc_clock_reset.reset_n
		.avs_hc_writedata_iDATA    (mm_interconnect_0_isp1362_if_0_hc_writedata),   //             hc.writedata
		.avs_hc_readdata_oDATA     (mm_interconnect_0_isp1362_if_0_hc_readdata),    //               .readdata
		.avs_hc_address_iADDR      (mm_interconnect_0_isp1362_if_0_hc_address),     //               .address
		.avs_hc_read_n_iRD_N       (~mm_interconnect_0_isp1362_if_0_hc_read),       //               .read_n
		.avs_hc_write_n_iWR_N      (~mm_interconnect_0_isp1362_if_0_hc_write),      //               .write_n
		.avs_hc_chipselect_n_iCS_N (~mm_interconnect_0_isp1362_if_0_hc_chipselect), //               .chipselect_n
		.avs_hc_irq_n_oINT0_N      (irq_mapper_receiver2_irq),                      //         hc_irq.irq_n
		.avs_dc_clk_iCLK           (altpll_sys),                                    //       dc_clock.clk
		.avs_dc_reset_n_iRST_N     (~rst_controller_reset_out_reset),               // dc_clock_reset.reset_n
		.avs_dc_writedata_iDATA    (mm_interconnect_0_isp1362_if_0_dc_writedata),   //             dc.writedata
		.avs_dc_readdata_oDATA     (mm_interconnect_0_isp1362_if_0_dc_readdata),    //               .readdata
		.avs_dc_address_iADDR      (mm_interconnect_0_isp1362_if_0_dc_address),     //               .address
		.avs_dc_read_n_iRD_N       (~mm_interconnect_0_isp1362_if_0_dc_read),       //               .read_n
		.avs_dc_write_n_iWR_N      (~mm_interconnect_0_isp1362_if_0_dc_write),      //               .write_n
		.avs_dc_chipselect_n_iCS_N (~mm_interconnect_0_isp1362_if_0_dc_chipselect), //               .chipselect_n
		.avs_dc_irq_n_oINT0_N      (irq_mapper_receiver1_irq),                      //         dc_irq.irq_n
		.USB_DATA                  (usb_conduit_end_DATA),                          //    conduit_end.export
		.USB_ADDR                  (usb_conduit_end_ADDR),                          //               .export
		.USB_RD_N                  (usb_conduit_end_RD_N),                          //               .export
		.USB_WR_N                  (usb_conduit_end_WR_N),                          //               .export
		.USB_CS_N                  (usb_conduit_end_CS_N),                          //               .export
		.USB_RST_N                 (usb_conduit_end_RST_N),                         //               .export
		.USB_INT0                  (usb_conduit_end_INT0),                          //               .export
		.USB_INT1                  (usb_conduit_end_INT1)                           //               .export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (22),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io (
		.m0_clk           (altpll_io),                                            //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                   // m0_reset.reset
		.s0_clk           (altpll_sys),                                           //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_m0_debugaccess)                      //         .debugaccess
	);

	DE2_115_SOPC_cpu cpu (
		.clk                                 (altpll_sys),                                        //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	DE2_115_SOPC_jtag_uart jtag_uart (
		.clk            (altpll_sys),                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver6_irq)                                   //               irq.irq
	);

	DE2_115_SOPC_key key (
		.clk        (altpll_io),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (in_port_to_the_key),                  // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)    //                 irq.irq
	);

	DE2_115_SOPC_lcd lcd (
		.reset_n       (~rst_controller_001_reset_out_reset),               //         reset.reset_n
		.clk           (altpll_io),                                         //           clk.clk
		.begintransfer (mm_interconnect_1_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_1_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_1_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_1_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_1_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_1_lcd_control_slave_address),       //              .address
		.LCD_RS        (LCD_RS_from_the_lcd),                               //      external.export
		.LCD_RW        (LCD_RW_from_the_lcd),                               //              .export
		.LCD_data      (LCD_data_to_and_from_the_lcd),                      //              .export
		.LCD_E         (LCD_E_from_the_lcd)                                 //              .export
	);

	DE2_115_SOPC_lcd_64_to_8_bits_dfa lcd_64_to_8_bits_dfa (
		.clk               (c3_out_clk_clk),                         //   clk.clk
		.reset_n           (~rst_controller_002_reset_out_reset),    // reset.reset_n
		.in_data           (lcd_ta_fifo_to_dfa_out_data),            //    in.data
		.in_valid          (lcd_ta_fifo_to_dfa_out_valid),           //      .valid
		.in_ready          (lcd_ta_fifo_to_dfa_out_ready),           //      .ready
		.in_startofpacket  (lcd_ta_fifo_to_dfa_out_startofpacket),   //      .startofpacket
		.in_endofpacket    (lcd_ta_fifo_to_dfa_out_endofpacket),     //      .endofpacket
		.in_empty          (lcd_ta_fifo_to_dfa_out_empty),           //      .empty
		.out_data          (lcd_64_to_8_bits_dfa_out_data),          //   out.data
		.out_valid         (lcd_64_to_8_bits_dfa_out_valid),         //      .valid
		.out_ready         (lcd_64_to_8_bits_dfa_out_ready),         //      .ready
		.out_startofpacket (lcd_64_to_8_bits_dfa_out_startofpacket), //      .startofpacket
		.out_endofpacket   (lcd_64_to_8_bits_dfa_out_endofpacket),   //      .endofpacket
		.out_empty         (lcd_64_to_8_bits_dfa_out_empty)          //      .empty
	);

	altera_avalon_pixel_converter #(
		.SOURCE_SYMBOLS_PER_BEAT (3)
	) lcd_pixel_converter (
		.clk       (c3_out_clk_clk),                         //       clk.clk
		.reset_n   (~rst_controller_002_reset_out_reset),    // clk_reset.reset_n
		.ready_out (lcd_64_to_8_bits_dfa_out_ready),         //        in.ready
		.valid_in  (lcd_64_to_8_bits_dfa_out_valid),         //          .valid
		.data_in   (lcd_64_to_8_bits_dfa_out_data),          //          .data
		.eop_in    (lcd_64_to_8_bits_dfa_out_endofpacket),   //          .endofpacket
		.sop_in    (lcd_64_to_8_bits_dfa_out_startofpacket), //          .startofpacket
		.empty_in  (lcd_64_to_8_bits_dfa_out_empty),         //          .empty
		.ready_in  (lcd_pixel_converter_out_ready),          //       out.ready
		.valid_out (lcd_pixel_converter_out_valid),          //          .valid
		.data_out  (lcd_pixel_converter_out_data),           //          .data
		.eop_out   (lcd_pixel_converter_out_endofpacket),    //          .endofpacket
		.sop_out   (lcd_pixel_converter_out_startofpacket),  //          .startofpacket
		.empty_out (lcd_pixel_converter_out_empty)           //          .empty
	);

	DE2_115_SOPC_lcd_pixel_fifo lcd_pixel_fifo (
		.wrclock                       (altpll_sys),                             //    clk_in.clk
		.wrreset_n                     (~rst_controller_reset_out_reset),        //  reset_in.reset_n
		.rdclock                       (c3_out_clk_clk),                         //   clk_out.clk
		.rdreset_n                     (~rst_controller_002_reset_out_reset),    // reset_out.reset_n
		.avalonst_sink_valid           (lcd_ta_sgdma_to_fifo_out_valid),         //        in.valid
		.avalonst_sink_data            (lcd_ta_sgdma_to_fifo_out_data),          //          .data
		.avalonst_sink_startofpacket   (lcd_ta_sgdma_to_fifo_out_startofpacket), //          .startofpacket
		.avalonst_sink_endofpacket     (lcd_ta_sgdma_to_fifo_out_endofpacket),   //          .endofpacket
		.avalonst_sink_empty           (lcd_ta_sgdma_to_fifo_out_empty),         //          .empty
		.avalonst_sink_ready           (lcd_ta_sgdma_to_fifo_out_ready),         //          .ready
		.avalonst_source_valid         (lcd_pixel_fifo_out_valid),               //       out.valid
		.avalonst_source_data          (lcd_pixel_fifo_out_data),                //          .data
		.avalonst_source_startofpacket (lcd_pixel_fifo_out_startofpacket),       //          .startofpacket
		.avalonst_source_endofpacket   (lcd_pixel_fifo_out_endofpacket),         //          .endofpacket
		.avalonst_source_empty         (lcd_pixel_fifo_out_empty),               //          .empty
		.avalonst_source_ready         (lcd_pixel_fifo_out_ready)                //          .ready
	);

	DE2_115_SOPC_lcd_sgdma lcd_sgdma (
		.clk                           (altpll_sys),                                 //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),            //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_lcd_sgdma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_lcd_sgdma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_lcd_sgdma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_lcd_sgdma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_lcd_sgdma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_lcd_sgdma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (lcd_sgdma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (lcd_sgdma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (lcd_sgdma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (lcd_sgdma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (lcd_sgdma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (lcd_sgdma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (lcd_sgdma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (lcd_sgdma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (lcd_sgdma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                   //          csr_irq.irq
		.m_read_readdata               (lcd_sgdma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (lcd_sgdma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (lcd_sgdma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (lcd_sgdma_m_read_address),                   //                 .address
		.m_read_read                   (lcd_sgdma_m_read_read),                      //                 .read
		.out_data                      (lcd_sgdma_out_data),                         //              out.data
		.out_valid                     (lcd_sgdma_out_valid),                        //                 .valid
		.out_ready                     (lcd_sgdma_out_ready),                        //                 .ready
		.out_endofpacket               (lcd_sgdma_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (lcd_sgdma_out_startofpacket),                //                 .startofpacket
		.out_empty                     (lcd_sgdma_out_empty)                         //                 .empty
	);

	DE2_115_SOPC_lcd_ta_fifo_to_dfa lcd_ta_fifo_to_dfa (
		.clk               (c3_out_clk_clk),                       //   clk.clk
		.reset_n           (~rst_controller_002_reset_out_reset),  // reset.reset_n
		.in_data           (lcd_pixel_fifo_out_data),              //    in.data
		.in_valid          (lcd_pixel_fifo_out_valid),             //      .valid
		.in_ready          (lcd_pixel_fifo_out_ready),             //      .ready
		.in_startofpacket  (lcd_pixel_fifo_out_startofpacket),     //      .startofpacket
		.in_endofpacket    (lcd_pixel_fifo_out_endofpacket),       //      .endofpacket
		.in_empty          (lcd_pixel_fifo_out_empty),             //      .empty
		.out_data          (lcd_ta_fifo_to_dfa_out_data),          //   out.data
		.out_valid         (lcd_ta_fifo_to_dfa_out_valid),         //      .valid
		.out_ready         (lcd_ta_fifo_to_dfa_out_ready),         //      .ready
		.out_startofpacket (lcd_ta_fifo_to_dfa_out_startofpacket), //      .startofpacket
		.out_endofpacket   (lcd_ta_fifo_to_dfa_out_endofpacket),   //      .endofpacket
		.out_empty         (lcd_ta_fifo_to_dfa_out_empty)          //      .empty
	);

	DE2_115_SOPC_lcd_ta_sgdma_to_fifo lcd_ta_sgdma_to_fifo (
		.clk               (altpll_sys),                                //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset),           // reset.reset_n
		.in_data           (avalon_st_adapter_001_out_0_data),          //    in.data
		.in_valid          (avalon_st_adapter_001_out_0_valid),         //      .valid
		.in_ready          (avalon_st_adapter_001_out_0_ready),         //      .ready
		.in_startofpacket  (avalon_st_adapter_001_out_0_startofpacket), //      .startofpacket
		.in_endofpacket    (avalon_st_adapter_001_out_0_endofpacket),   //      .endofpacket
		.in_empty          (avalon_st_adapter_001_out_0_empty),         //      .empty
		.out_data          (lcd_ta_sgdma_to_fifo_out_data),             //   out.data
		.out_valid         (lcd_ta_sgdma_to_fifo_out_valid),            //      .valid
		.out_ready         (lcd_ta_sgdma_to_fifo_out_ready),            //      .ready
		.out_startofpacket (lcd_ta_sgdma_to_fifo_out_startofpacket),    //      .startofpacket
		.out_endofpacket   (lcd_ta_sgdma_to_fifo_out_endofpacket),      //      .endofpacket
		.out_empty         (lcd_ta_sgdma_to_fifo_out_empty)             //      .empty
	);

	DE2_115_SOPC_ledg ledg (
		.clk        (altpll_io),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledg_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_ledg)                // external_connection.export
	);

	DE2_115_SOPC_ledr ledr (
		.clk        (altpll_io),                            //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_1_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ledr_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_ledr)                // external_connection.export
	);

	DE2_115_SOPC_pll pll (
		.clk                (clk_50),                                    //       inclk_interface.clk
		.reset              (rst_controller_003_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_sys),                                //                    c0.clk
		.c1                 (altpll_sdram),                              //                    c1.clk
		.c2                 (altpll_io),                                 //                    c2.clk
		.c3                 (c3_out_clk_clk),                            //                    c3.clk
		.areset             (pll_areset_conduit_export),                 //        areset_conduit.export
		.locked             (locked_from_the_pll),                       //        locked_conduit.export
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.phasedone          (),                                          //           (terminated)
		.phasecounterselect (4'b0000),                                   //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0)                                       //           (terminated)
	);

	DE2_115_SOPC_sdram sdram (
		.clk            (altpll_sys),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	SEG7_IF #(
		.SEG7_NUM       (8),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.s_address   (mm_interconnect_1_seg7_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_1_seg7_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_1_seg7_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_1_seg7_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_1_seg7_avalon_slave_writedata), //                 .writedata
		.SEG7        (SEG7_from_the_seg7),                            //      conduit_end.export
		.s_clk       (altpll_io),                                     //       clock_sink.clk
		.s_reset     (rst_controller_001_reset_out_reset)             // clock_sink_reset.reset
	);

	DE2_115_SOPC_sw sw (
		.clk        (altpll_io),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port    (in_port_to_the_sw),                   // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)    //                 irq.irq
	);

	DE2_115_SOPC_sysid sysid (
		.clock    (altpll_io),                                      //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DE2_115_SOPC_timer timer (
		.clk        (altpll_io),                             //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)          //   irq.irq
	);

	DE2_115_SOPC_timer_stamp timer_stamp (
		.clk        (altpll_sys),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             // reset.reset_n
		.address    (mm_interconnect_0_timer_stamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_stamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_stamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_stamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_stamp_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver7_irq)                     //   irq.irq
	);

	DE2_115_SOPC_vga vga (
		.clk           (c3_out_clk_clk),                                        //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                    //              reset.reset
		.data          (video_rgb_resampler_0_avalon_rgb_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                   .endofpacket
		.valid         (video_rgb_resampler_0_avalon_rgb_source_valid),         //                   .valid
		.ready         (video_rgb_resampler_0_avalon_rgb_source_ready),         //                   .ready
		.VGA_CLK       (vga_data_CLK),                                          // external_interface.export
		.VGA_HS        (vga_data_HS),                                           //                   .export
		.VGA_VS        (vga_data_VS),                                           //                   .export
		.VGA_BLANK     (vga_data_BLANK),                                        //                   .export
		.VGA_SYNC      (vga_data_SYNC),                                         //                   .export
		.VGA_R         (vga_data_R),                                            //                   .export
		.VGA_G         (vga_data_G),                                            //                   .export
		.VGA_B         (vga_data_B)                                             //                   .export
	);

	DE2_115_SOPC_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (c3_out_clk_clk),                                        //               clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                    //             reset.reset
		.stream_in_startofpacket  (avalon_st_adapter_out_0_startofpacket),                 //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (avalon_st_adapter_out_0_endofpacket),                   //                  .endofpacket
		.stream_in_valid          (avalon_st_adapter_out_0_valid),                         //                  .valid
		.stream_in_ready          (avalon_st_adapter_out_0_ready),                         //                  .ready
		.stream_in_data           (avalon_st_adapter_out_0_data),                          //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)           //                  .data
	);

	DE2_115_SOPC_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                        (clk_50),                                                    //                                      clk_50_clk.clk
		.pll_c0_clk                                            (altpll_sys),                                                //                                          pll_c0.clk
		.pll_c2_clk                                            (altpll_io),                                                 //                                          pll_c2.clk
		.cpu_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                            //                 cpu_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                        // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.timer_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                        //               timer_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                               (cpu_data_master_address),                                   //                                 cpu_data_master.address
		.cpu_data_master_waitrequest                           (cpu_data_master_waitrequest),                               //                                                .waitrequest
		.cpu_data_master_byteenable                            (cpu_data_master_byteenable),                                //                                                .byteenable
		.cpu_data_master_read                                  (cpu_data_master_read),                                      //                                                .read
		.cpu_data_master_readdata                              (cpu_data_master_readdata),                                  //                                                .readdata
		.cpu_data_master_readdatavalid                         (cpu_data_master_readdatavalid),                             //                                                .readdatavalid
		.cpu_data_master_write                                 (cpu_data_master_write),                                     //                                                .write
		.cpu_data_master_writedata                             (cpu_data_master_writedata),                                 //                                                .writedata
		.cpu_data_master_debugaccess                           (cpu_data_master_debugaccess),                               //                                                .debugaccess
		.cpu_instruction_master_address                        (cpu_instruction_master_address),                            //                          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                        //                                                .waitrequest
		.cpu_instruction_master_read                           (cpu_instruction_master_read),                               //                                                .read
		.cpu_instruction_master_readdata                       (cpu_instruction_master_readdata),                           //                                                .readdata
		.cpu_instruction_master_readdatavalid                  (cpu_instruction_master_readdatavalid),                      //                                                .readdatavalid
		.lcd_sgdma_descriptor_read_address                     (lcd_sgdma_descriptor_read_address),                         //                       lcd_sgdma_descriptor_read.address
		.lcd_sgdma_descriptor_read_waitrequest                 (lcd_sgdma_descriptor_read_waitrequest),                     //                                                .waitrequest
		.lcd_sgdma_descriptor_read_read                        (lcd_sgdma_descriptor_read_read),                            //                                                .read
		.lcd_sgdma_descriptor_read_readdata                    (lcd_sgdma_descriptor_read_readdata),                        //                                                .readdata
		.lcd_sgdma_descriptor_read_readdatavalid               (lcd_sgdma_descriptor_read_readdatavalid),                   //                                                .readdatavalid
		.lcd_sgdma_descriptor_write_address                    (lcd_sgdma_descriptor_write_address),                        //                      lcd_sgdma_descriptor_write.address
		.lcd_sgdma_descriptor_write_waitrequest                (lcd_sgdma_descriptor_write_waitrequest),                    //                                                .waitrequest
		.lcd_sgdma_descriptor_write_write                      (lcd_sgdma_descriptor_write_write),                          //                                                .write
		.lcd_sgdma_descriptor_write_writedata                  (lcd_sgdma_descriptor_write_writedata),                      //                                                .writedata
		.lcd_sgdma_m_read_address                              (lcd_sgdma_m_read_address),                                  //                                lcd_sgdma_m_read.address
		.lcd_sgdma_m_read_waitrequest                          (lcd_sgdma_m_read_waitrequest),                              //                                                .waitrequest
		.lcd_sgdma_m_read_read                                 (lcd_sgdma_m_read_read),                                     //                                                .read
		.lcd_sgdma_m_read_readdata                             (lcd_sgdma_m_read_readdata),                                 //                                                .readdata
		.lcd_sgdma_m_read_readdatavalid                        (lcd_sgdma_m_read_readdatavalid),                            //                                                .readdatavalid
		.clock_crossing_io_s0_address                          (mm_interconnect_0_clock_crossing_io_s0_address),            //                            clock_crossing_io_s0.address
		.clock_crossing_io_s0_write                            (mm_interconnect_0_clock_crossing_io_s0_write),              //                                                .write
		.clock_crossing_io_s0_read                             (mm_interconnect_0_clock_crossing_io_s0_read),               //                                                .read
		.clock_crossing_io_s0_readdata                         (mm_interconnect_0_clock_crossing_io_s0_readdata),           //                                                .readdata
		.clock_crossing_io_s0_writedata                        (mm_interconnect_0_clock_crossing_io_s0_writedata),          //                                                .writedata
		.clock_crossing_io_s0_burstcount                       (mm_interconnect_0_clock_crossing_io_s0_burstcount),         //                                                .burstcount
		.clock_crossing_io_s0_byteenable                       (mm_interconnect_0_clock_crossing_io_s0_byteenable),         //                                                .byteenable
		.clock_crossing_io_s0_readdatavalid                    (mm_interconnect_0_clock_crossing_io_s0_readdatavalid),      //                                                .readdatavalid
		.clock_crossing_io_s0_waitrequest                      (mm_interconnect_0_clock_crossing_io_s0_waitrequest),        //                                                .waitrequest
		.clock_crossing_io_s0_debugaccess                      (mm_interconnect_0_clock_crossing_io_s0_debugaccess),        //                                                .debugaccess
		.cpu_debug_mem_slave_address                           (mm_interconnect_0_cpu_debug_mem_slave_address),             //                             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                             (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                                .write
		.cpu_debug_mem_slave_read                              (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                                .read
		.cpu_debug_mem_slave_readdata                          (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                                .readdata
		.cpu_debug_mem_slave_writedata                         (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                                .writedata
		.cpu_debug_mem_slave_byteenable                        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                                .byteenable
		.cpu_debug_mem_slave_waitrequest                       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                                .waitrequest
		.cpu_debug_mem_slave_debugaccess                       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                                .debugaccess
		.ISP1362_IF_0_dc_address                               (mm_interconnect_0_isp1362_if_0_dc_address),                 //                                 ISP1362_IF_0_dc.address
		.ISP1362_IF_0_dc_write                                 (mm_interconnect_0_isp1362_if_0_dc_write),                   //                                                .write
		.ISP1362_IF_0_dc_read                                  (mm_interconnect_0_isp1362_if_0_dc_read),                    //                                                .read
		.ISP1362_IF_0_dc_readdata                              (mm_interconnect_0_isp1362_if_0_dc_readdata),                //                                                .readdata
		.ISP1362_IF_0_dc_writedata                             (mm_interconnect_0_isp1362_if_0_dc_writedata),               //                                                .writedata
		.ISP1362_IF_0_dc_chipselect                            (mm_interconnect_0_isp1362_if_0_dc_chipselect),              //                                                .chipselect
		.ISP1362_IF_0_hc_address                               (mm_interconnect_0_isp1362_if_0_hc_address),                 //                                 ISP1362_IF_0_hc.address
		.ISP1362_IF_0_hc_write                                 (mm_interconnect_0_isp1362_if_0_hc_write),                   //                                                .write
		.ISP1362_IF_0_hc_read                                  (mm_interconnect_0_isp1362_if_0_hc_read),                    //                                                .read
		.ISP1362_IF_0_hc_readdata                              (mm_interconnect_0_isp1362_if_0_hc_readdata),                //                                                .readdata
		.ISP1362_IF_0_hc_writedata                             (mm_interconnect_0_isp1362_if_0_hc_writedata),               //                                                .writedata
		.ISP1362_IF_0_hc_chipselect                            (mm_interconnect_0_isp1362_if_0_hc_chipselect),              //                                                .chipselect
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.lcd_sgdma_csr_address                                 (mm_interconnect_0_lcd_sgdma_csr_address),                   //                                   lcd_sgdma_csr.address
		.lcd_sgdma_csr_write                                   (mm_interconnect_0_lcd_sgdma_csr_write),                     //                                                .write
		.lcd_sgdma_csr_read                                    (mm_interconnect_0_lcd_sgdma_csr_read),                      //                                                .read
		.lcd_sgdma_csr_readdata                                (mm_interconnect_0_lcd_sgdma_csr_readdata),                  //                                                .readdata
		.lcd_sgdma_csr_writedata                               (mm_interconnect_0_lcd_sgdma_csr_writedata),                 //                                                .writedata
		.lcd_sgdma_csr_chipselect                              (mm_interconnect_0_lcd_sgdma_csr_chipselect),                //                                                .chipselect
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                   //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                     //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                      //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                  //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                 //                                                .writedata
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                        //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                          //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                           //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                       //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                      //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                     //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                    //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect),                     //                                                .chipselect
		.timer_s1_address                                      (mm_interconnect_0_timer_s1_address),                        //                                        timer_s1.address
		.timer_s1_write                                        (mm_interconnect_0_timer_s1_write),                          //                                                .write
		.timer_s1_readdata                                     (mm_interconnect_0_timer_s1_readdata),                       //                                                .readdata
		.timer_s1_writedata                                    (mm_interconnect_0_timer_s1_writedata),                      //                                                .writedata
		.timer_s1_chipselect                                   (mm_interconnect_0_timer_s1_chipselect),                     //                                                .chipselect
		.timer_stamp_s1_address                                (mm_interconnect_0_timer_stamp_s1_address),                  //                                  timer_stamp_s1.address
		.timer_stamp_s1_write                                  (mm_interconnect_0_timer_stamp_s1_write),                    //                                                .write
		.timer_stamp_s1_readdata                               (mm_interconnect_0_timer_stamp_s1_readdata),                 //                                                .readdata
		.timer_stamp_s1_writedata                              (mm_interconnect_0_timer_stamp_s1_writedata),                //                                                .writedata
		.timer_stamp_s1_chipselect                             (mm_interconnect_0_timer_stamp_s1_chipselect)                //                                                .chipselect
	);

	DE2_115_SOPC_mm_interconnect_1 mm_interconnect_1 (
		.pll_c2_clk                                             (altpll_io),                                         //                                           pll_c2.clk
		.clock_crossing_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                // clock_crossing_io_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_m0_address                           (clock_crossing_io_m0_address),                      //                             clock_crossing_io_m0.address
		.clock_crossing_io_m0_waitrequest                       (clock_crossing_io_m0_waitrequest),                  //                                                 .waitrequest
		.clock_crossing_io_m0_burstcount                        (clock_crossing_io_m0_burstcount),                   //                                                 .burstcount
		.clock_crossing_io_m0_byteenable                        (clock_crossing_io_m0_byteenable),                   //                                                 .byteenable
		.clock_crossing_io_m0_read                              (clock_crossing_io_m0_read),                         //                                                 .read
		.clock_crossing_io_m0_readdata                          (clock_crossing_io_m0_readdata),                     //                                                 .readdata
		.clock_crossing_io_m0_readdatavalid                     (clock_crossing_io_m0_readdatavalid),                //                                                 .readdatavalid
		.clock_crossing_io_m0_write                             (clock_crossing_io_m0_write),                        //                                                 .write
		.clock_crossing_io_m0_writedata                         (clock_crossing_io_m0_writedata),                    //                                                 .writedata
		.clock_crossing_io_m0_debugaccess                       (clock_crossing_io_m0_debugaccess),                  //                                                 .debugaccess
		.key_s1_address                                         (mm_interconnect_1_key_s1_address),                  //                                           key_s1.address
		.key_s1_write                                           (mm_interconnect_1_key_s1_write),                    //                                                 .write
		.key_s1_readdata                                        (mm_interconnect_1_key_s1_readdata),                 //                                                 .readdata
		.key_s1_writedata                                       (mm_interconnect_1_key_s1_writedata),                //                                                 .writedata
		.key_s1_chipselect                                      (mm_interconnect_1_key_s1_chipselect),               //                                                 .chipselect
		.lcd_control_slave_address                              (mm_interconnect_1_lcd_control_slave_address),       //                                lcd_control_slave.address
		.lcd_control_slave_write                                (mm_interconnect_1_lcd_control_slave_write),         //                                                 .write
		.lcd_control_slave_read                                 (mm_interconnect_1_lcd_control_slave_read),          //                                                 .read
		.lcd_control_slave_readdata                             (mm_interconnect_1_lcd_control_slave_readdata),      //                                                 .readdata
		.lcd_control_slave_writedata                            (mm_interconnect_1_lcd_control_slave_writedata),     //                                                 .writedata
		.lcd_control_slave_begintransfer                        (mm_interconnect_1_lcd_control_slave_begintransfer), //                                                 .begintransfer
		.ledg_s1_address                                        (mm_interconnect_1_ledg_s1_address),                 //                                          ledg_s1.address
		.ledg_s1_write                                          (mm_interconnect_1_ledg_s1_write),                   //                                                 .write
		.ledg_s1_readdata                                       (mm_interconnect_1_ledg_s1_readdata),                //                                                 .readdata
		.ledg_s1_writedata                                      (mm_interconnect_1_ledg_s1_writedata),               //                                                 .writedata
		.ledg_s1_chipselect                                     (mm_interconnect_1_ledg_s1_chipselect),              //                                                 .chipselect
		.ledr_s1_address                                        (mm_interconnect_1_ledr_s1_address),                 //                                          ledr_s1.address
		.ledr_s1_write                                          (mm_interconnect_1_ledr_s1_write),                   //                                                 .write
		.ledr_s1_readdata                                       (mm_interconnect_1_ledr_s1_readdata),                //                                                 .readdata
		.ledr_s1_writedata                                      (mm_interconnect_1_ledr_s1_writedata),               //                                                 .writedata
		.ledr_s1_chipselect                                     (mm_interconnect_1_ledr_s1_chipselect),              //                                                 .chipselect
		.seg7_avalon_slave_address                              (mm_interconnect_1_seg7_avalon_slave_address),       //                                seg7_avalon_slave.address
		.seg7_avalon_slave_write                                (mm_interconnect_1_seg7_avalon_slave_write),         //                                                 .write
		.seg7_avalon_slave_read                                 (mm_interconnect_1_seg7_avalon_slave_read),          //                                                 .read
		.seg7_avalon_slave_readdata                             (mm_interconnect_1_seg7_avalon_slave_readdata),      //                                                 .readdata
		.seg7_avalon_slave_writedata                            (mm_interconnect_1_seg7_avalon_slave_writedata),     //                                                 .writedata
		.sw_s1_address                                          (mm_interconnect_1_sw_s1_address),                   //                                            sw_s1.address
		.sw_s1_write                                            (mm_interconnect_1_sw_s1_write),                     //                                                 .write
		.sw_s1_readdata                                         (mm_interconnect_1_sw_s1_readdata),                  //                                                 .readdata
		.sw_s1_writedata                                        (mm_interconnect_1_sw_s1_writedata),                 //                                                 .writedata
		.sw_s1_chipselect                                       (mm_interconnect_1_sw_s1_chipselect),                //                                                 .chipselect
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),     //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata)     //                                                 .readdata
	);

	DE2_115_SOPC_irq_mapper irq_mapper (
		.clk           (altpll_sys),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (~irq_mapper_receiver1_irq),      // receiver1.irq
		.receiver2_irq (~irq_mapper_receiver2_irq),      // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_io),                          //       receiver_clk.clk
		.sender_clk     (altpll_sys),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	DE2_115_SOPC_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (c3_out_clk_clk),                        // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_002_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (lcd_pixel_converter_out_data),          //     in_0.data
		.in_0_valid          (lcd_pixel_converter_out_valid),         //         .valid
		.in_0_ready          (lcd_pixel_converter_out_ready),         //         .ready
		.in_0_startofpacket  (lcd_pixel_converter_out_startofpacket), //         .startofpacket
		.in_0_endofpacket    (lcd_pixel_converter_out_endofpacket),   //         .endofpacket
		.in_0_empty          (lcd_pixel_converter_out_empty),         //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)    //         .endofpacket
	);

	DE2_115_SOPC_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (altpll_sys),                                // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (lcd_sgdma_out_data),                        //     in_0.data
		.in_0_valid          (lcd_sgdma_out_valid),                       //         .valid
		.in_0_ready          (lcd_sgdma_out_ready),                       //         .ready
		.in_0_startofpacket  (lcd_sgdma_out_startofpacket),               //         .startofpacket
		.in_0_endofpacket    (lcd_sgdma_out_endofpacket),                 //         .endofpacket
		.in_0_empty          (lcd_sgdma_out_empty),                       //         .empty
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)          //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_sys),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (altpll_io),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (c3_out_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
